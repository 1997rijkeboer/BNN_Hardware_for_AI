-- Top-level testbench
-- Loads in constant weights, others from TCL script

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity top_tb is
    generic (
        INPUT_WIDTH     : integer := 8;
        OUTPUT_WIDTH    : integer := 4;
        INPUT_COLS      : integer := 28;
        INPUT_ROWS      : integer := 28;
        OUTPUT_COLS     : integer := 1
    );
    port (
        -- System
        reset       : in  std_logic;

        -- Input data
        row_in      : in  std_logic_vector(INPUT_COLS*INPUT_WIDTH-1 downto 0);
        ready       : in  std_logic;

        -- Output data
        row_out     : out std_logic_vector(OUTPUT_COLS*OUTPUT_WIDTH-1 downto 0);
        done        : out std_logic
    );
end entity;


architecture sim of top_tb is

    constant CLK_PERIOD : time := 10 ns;

    signal clk : std_logic := '0';

    signal w_en, w_in, w_out : std_logic;

    constant WEIGHTS : std_logic_vector(0 to 49362-1) := "001001000010111110000111111010111110111000000110110110001010010000011111101101000011111111001110010001111110001111111101000001010011111111111110110111100001011111110111110101100000110111110010111111111111100100000100010111111101000010100100001111011110010111111001110100000010110001001001100100000010111000011111010111011001010111111111101001111110100010111111111111111010110110000000000001011111000011101011011111100000000001110100000000000001111101000000000011011111100010000011011111001011111010000000011011111011001100001001110001011110011011111000000000000001110011011111000000010000000000001111111100010000000000000000000001001111101000000000001111100110010010010000000000011111001011111011001111001111110000000000001000000001111110001011111111111111000000000111111001000000000111111001000000000000000000000000000111010000000000000111111000000000000111011011111111000000000000111111000111101010111111011111111010111111001000000000001001000111111001110111110000000000111111011000000000000000000000100000101110011011001000000001000000000000000000000000000000100111011000111110111111010000000000110110110111110000111111011000000000000000000100110111100101011100100111000000100100100001000000000000010111000000000100000111000000100100000111100110111001000100100000111100000011000110011010111011100100111000000000100000011100111111101000010100100000100111111001000100000001000101000100100111111000000000100100000010000000000000100100000000100110010000000110100100111001000100101101110100110111000000111000000000010110010000001000000011000000001001010010000000001000010000100001011011000100100000001001110110110000001011000000001011001000001011001100001001000000001000011011000001001010000100000000000000001001000000000110100001001001001010100010010010000000000000000001001000000000110111110010100110010100010010010001000001001000000011000000001000000000000000010001001001000001001000011000000000000101001111001001011111011111000000000111011011000000000001011100100000000101011111000000000101011111111011111000000000001001110101001111111011111111011111111001111000000000000001011101001111001000000100000000101011111000000000000000000000000000111011111000000000000000010000000000000000000100001011111001101110111101111011100000000000110101101001011110101001100000000000010000110001111011011001111111111011010000100101111110010000000011111011000000100011111001000000101011111111011111011010000100011111011001111001101111111011111111101111111000000111001000011011111111101101101100000101111111111010000100010000000000000101111111111100000000001111011110000100010000100000011001011111011001001101011111011010000000001111101011001011001111001000100000000000000000000000000000000100100011000000000000000000000000000000100001000000000100000100111110111100000000100010011000000000000101000111111111011100000001100001100100000000000000000000000100110000111111111000001011100100000000000000000000000111111111000110011000000000000000000000000110000000000000000000000000000111111111100110000000000000111111111100100000111111111000000000010000010011011110011111110011010110000000010101010100110000010111110111000000010011111111000100100011110110011111111010000010011110110001010110011011110011110111011111111100000010011010110011110110001001111000001000011111110100000000000100000001000110011111110011100000011111111000000010000000000011110110011011111011001110011111111100000010001011010011111110011010111111111100001101101110010000000000000110010000011101001000000100010001100100000000111001111110010000010110010110000000110010000001100111010010000110010000110010000100010000110010000101001101010000000110010000010100011011011111010010000011101101011101001110110000010010000000000000010000101111100110011001101100000000010010000110111000110000000111101010110111000010010000110000000010001100100100111001001011000001011001001001100110101000001011111110000001001011110100111001000011100000000001000001001001011110110111001001010001001001001001001001001110000001001100100000000001011001001011010000000100110010001001010100100001110110111000000000000001001111110111100000000100010110100110101001011010000001001000000000001011011000000001000000101001001000001001001100011001000000000111011100000000000111001100000010000000000000000000000111011000000000000111011000111001100111011000111001000000000000011001000111001000111001000111001000111001000000001000000000000111001000111111111011110011111001000000100001001001101100111111111001000000011000111110110000000000000000000000000000111001000110111001111001000000100000110111111101001100111001000000000000001000000111011001110011011111011111000000000110011011000001000110100011001000000110010001001000000110110001110110011001100110110111011110111011110110011110110011111110011001000000100000011110000011011101000101100000110011001000000000001001000000001000111011001001000000111011000000000000000000000000000011110000011100000101110010011000000000100101010110011001110110001100001000001000000110010110010000110110010001101011100000000010000000000100100111000000000110000100000000100110100100110110100000000000110100111100000000110000010000100110110010100000000000110010100110100101010010000000000000110100111001011001000000000110000100010110110000000000000000000100001000001001000010010010110110110110000000110000111000000000110100001110100101110000100000010110000000000000000000000101111000010100010000000000000000000000010000000000100010010000000100000000000000000000000000000110000000000100100000000100000000000000100000000010100000001000000000000000110000010010110110011000000000000101100000000011000000000100000100001110011000000000000000000000101100000000001011000000000000000110000110000100000110000100110000100110000000100000000000000000000001101001000001000001001011010000000101001011000000000001011101000000000001001001001100100001011011001011101011000000001001101001101001001101001011011011001001001000000000001001001001001001000000000010000000001001001011000000000000001001000000101001001000000000000001001001000000010000001001011001001101001001001000001001101001000000000000000001001001001001001000000000000000100000111000001111000000111000001010000000101000000000000001111000000000100000111000000010000000111110000111001100000000001111000000111000000111000001111001000111000010000110000010000001111000000010111000000110001111000000000000111000100000000111001111000101000111111010000000000010000000000000010100000111010000001111001111000000000011000011001001111000000011001001100000000000000111111111111111111111111111000000000111111111000000000111111111000000000111111111000000000111111111111111111000000000111111111100000000111111111111111111111111111000000000111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000111111111000000000000000000111111111111111111000000000111111111000000000000000000111111111111111111111111111111110110001011011000111011001001001111010111011011011111110111011011011111110111001001001111010111000011011001001011111111111001011011000000011000001011001011011001001001111110111111111111001011011100000000100000000001011011111110111110110110000000100001011011111110101101111011111110110111110111011011111001001011000000001000001011010010110000000001001011011001001001111111111000001100111111111110111011111111011000001000111110001000001000111110011000001000111111010101101000111111011111111010000000100110100111111110101111110101111110011111111111000000100111110111111111011101000100101111100111111111000001000000001001100100100110111011000011000111110001001001100000000000111110010111111111111110111111110011000001010111100111110101011111111011111001001000000000000000111100001111000000111000000100000001111000001000000001111010011100001000111011001100001000111001001111010000000101001111000100111000001111001000111000100111000000000000000111001001111000010000000000000000001111010000100000000000000000000010001111000000000000000001010001000010000000000001100001101111011010001000001111001000100001010001000000111000000111000000000000000000001001001011010001001001001110000000011001011000000000001011010000000000001001011100001000001001011001001011000000000001011011001001001100001011011010010001001001000000000001001011001001011101101000000101100111011011100000000000000000000001000001001001000000000011011101010000000000000100001000001001001001000011010011001011000000000000001000111011011001001001110000001110110100011001011011011101011001011110110110000000111110111110001011011110110100011011111110110110011011111011010011110110110011011011011011011011001111011011111011001011110110110111000111001011111111001101010100011001011011110110110010110110111111111001011011100111110010000101110110110110110100001100111001000011011010111001011111110111111011011111001011111011001111000100000101001111000000000000000000000000000100011111001000000100000111001000000001010000000000010011010111000000000000000000100010110000000000001000000001000000001000000000000000100000111100000000000000000011010100001001001000000000100011111000000000000001000000000000001000000000000000000000000110011111000000000100100000000011011001000000000001001000011010000000000000000000011010000000001000111100000011000010111000000000001000011000000000011000111001001000001000111000000010010011111001000111000000000000000111000001111000000111000000111000001111000000000011000011000000111000000010111000000001110111000100000001000000000000110111000011000000000001000110000000000000100000001000101000000111001000111011000111000000000011000001011000111000000111000000110110111001000000100111111100011111100111111001001000110011111000000000100111111000000000100001111000000000100101111000011111001000000100111111110111111110110111100111111100110111001000000111011111000111111000000000111100000100111111001000000001000000000000000100111111110000100000000000000000000001001000111111111110111111100000111100011111000000000110100111100111111100101111000000000001000000100100100100101100000110100001000000100000100001000010100001001010000010110110100000000000100100100110110100000000000110110100010100100010100100110000000110100100010000000110111100110100100100110000000000000100110100001000000000000000010010000100111100000000000000000000000000010001000000000000100100100100010010001110110100000000000110100000110100100110110100000000000000110000111000000001010011111000000000000000101001011000110000111000010000100000111000000000000000111000000111000000000000000011000010111000000111000000111000000111000010000110000111010000111000000011001000000010101001000000000000000000100100011011100001000010000100000000000000100111110000000000100000000111000000111110010111010000000000000011011001001000010111000000000000000000000000010010110100101101110011111000000000000110000000000000010011100000000000111111101010000000110011101110011101000000000110111101101111100110110100010011101000010111000000000101111101110111101101000000000000000111110001000000000000000000111000001111011011000000000010000000000000000010000000000000000010010000001000001110111101111000000000000011111011101011111101100100000001001001110110110100010110110110110000000001110000110011010000100100111000000000110100110000000010110110110110110110000001001100100110111110010111110010100100110110110110000011001110110010110100110111011110001011011110010110000000000001000010000100100110010111000011000110011010000000000000000001110000001110010010111100110100110110000000000111100011110010110110100110010011010000000100011000010000011000011000010000000101001011010000001001010110110100000001011010010000000101011010010011010010000100001011010110001000010011011010010010110001001010000100001000000000001010010011000110000011010001010010000100000000000101010000100001001010000000001011010000000000101000000101000001011011001010001000010000010010101000001001000010011010010011010010101011110000000000111111111111111111111111111000000000111111111000000000000000000000000000000000000000000000000000000111111111111111111000000000111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000111010011000000000000000000000000000111110011000000000011010011000000000111111111000000000111111011000000000000000000111111111000000000000000000000000000000000000000000000111111011000000000000000000111110011111101101000000000111111111111111111111111011000000000111101111000000000111111011011111111000000000000000000110101011000000000011110111111111011110111111000000000101001100001111010000010000000010101000010011011000000000111101011000000000111011000000000000100011111000010000000011000011011001001000000010011000110000000110000000111011000000111101000000000000010000010011000000000100110101000010001001001000010111000000000000000000001111000000111110110111001000001010000111111011110110011000000000000110011000000000000000000000010101000100011001010100000000011111100000111000100111100000000001001110000000000000001111000000000000010111100001000000000111000100111000101000000000111000100111110100111110100111000100111100000000000001101000000111000000011100000010110100111000100000000001000000001000001001111000000000010111000000000000000000000000001100100000111100000111111001111000000000000011111101000111000000111100101000000000111111110000000000000000000000000000111111110000000000111111110000000000110111110000000000111111111000000000000000000011111111000000000000000000000000000000000000000000000111111110000000000000000000101101101111111111000000000111111110101111111111111111000000000111111111000000000111111110111111110000000000000000000000000000000000000111111111111101111000000000000000000000000000000001000111111001110111001111111001000000100111011001000001001111110011000000100111111011000000000111111010111111010100000010111100011111111011111111001111110011111100001111001111111111001111110011001110001001010000111111001000000100100001000001010000111111011000011101111001011100000000000000100111011111101111001011111111111110011000000100111111111111110011111111011110000000000000000010110000000100100010100101000000000000000100000000000110101001000000000110100111000000000010100101110100101000000000100100001010100000010100100010101001110110100000000000000000000110100011010001010010000000010101101000000000000000000011000000110110101000001000100110000000000000000000000000100000110110001011010011010110011010000000001000001010100001110100111000100000000000000111111011111011110111111111010000000111111111000010010110111011000000110111111101100000000111111011111111011001000010111111011111111111111111111111111011111111111000000010111111011111111011100000000011000000111111011001000000010000110100000000111111011000000100111111011000000000000000000111111111111111111100100000111111011000000110100000100111111011111111111010000000000000000011100000111100101011110000000000011111000101000000000111010001000000000011100000010010001011100000111110000101000011011000000111110100111110100111110001111110000000011001111110000011100000000101000000000000011000000000000000001000010000110010111100000000010001011010000000000000000000001011011000011110100001111000111100000101100101011111100011000100011110000000010010001000000010010000000000001000000000000000001000000000000000000000000001000000001000100000111011111000000000000000001001000001000000001111110110000000000000000001000000000000000000000000000000000001000000000111000000000000000000000001000000001000000000000000000000000000000000000000000001000000001000100000000100000110100010000000001110100100010000010000000001110110000000000000000000000111011011101000001011011011000000000001000001000000000110110011000000000011010011000000000111010001111010001000101001011010011111010111111011011110100011011000011000100000100000000011010011011111110000100000011010111000000000000100000000010100011011111000000000000010010000100000000000000100010011111001001010000000011000011000000000000000000011000011111010111100100111000000000011111111010101000011101110000000000000100100000000000111111101000000000011110101001000101011101101011110111000000000011110101011110110011110111111111101011101100000000000010100000111101101111111111000000100011111100000000000000100111111111101011101111100000110000100100100000000000000000000000000111101111111011111011111101100101001011111111111101101011110100000100100000001000101111111100111111101111111000000000100110111000001000100111111010000000101101111100000001100101111100111111000000000111111111111110111110101111100111110100111111000000000100100010101111111110000000111101011111111111000000000010001000111000000111111111000000000100000111000001001000000000100101110101111111101001111101111111000000000111101101100111111101101111000100011110100000011011111011111110011011111110100011011111110100000000011111111100100000011011111100100001011011111011011111100100000011011100001011111001011110011111111011011111100000000111111111011111111101001101000000001011111111110110010000000000001001011011111111000000000011111110110110111110100010001011110011011111001011011011111111100000000000000001011111111011011011111111111000000000100100000111110110101100010000000100110000110000000000111101011000000000101101000000000000101101000111101011000000000111101101101100000111100000111011011101110010000000000100110110111100000000000000000000000111100101000000000000000000000000000000000000000000000000000000000000000000000100101010000111100111000000000110100000000000000000000000111101000101100001000000000100101100000000000000000000000000000110111111000100000111110100000000000111110000000000000000101010000000000000000000111111111000000000000000000000000000000000000000000000110100100000000000000000000000001010110110100000000000110100111110010100000001000000000000110100100000000000010011111110110111110000000000000000000000000000000000110100100100100101000000000000000000000100000000000000111111111111111111111111111000000000111111111000000000111111111000000000111111111000000000111111111111111111000000000111111111111111111111111111111111111111111111000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111000000000111111111000000000000000000111111111111111111111111111111011011000000100000000001000000000101101111000000010111111011000000000001111011100000000111111110000000000000000000101111011000000000111100100000000000000000001000000100101011011000000000000000000111111110011111110000000100101101011101000111111111100000000100111111011000110000101001011101001111000000000000100100111110100000000000111111011111100100000000000111100100000000000000000000100100111000100111110100111000011000000100111000001000100000111000001000110100001000011000100100111110100111000000000100100111100100110100100110100000111110100110000001000000000110100100111110100000000000000100110111001001000000111000100100000100110111000011010000000000001001000001001100000110111100100100100000100100100111000000000100100000110100111100100000000010000000000001000000000000000000000000000100011001000000000010001000000000000010101001000000000000011001000000000000000000000000001000000100000000000100000000000000000000000000110001000000000000000000000101011001100001001000000000100001001001111101111011001000000000010011011000000000011001001100001001000000000000000000101001011000000000010001000100101111000000000000000000000000000000000000000100111000000011000001111011000000101011111000000000000110110000000000000100110000000000000100110000101111000000000011111110000010111001111111000110110000110111000000010000110111000111110110000000000000000011111110010000000000000000000000000001111111000000010000000000000010000010000000000111011010001110010001110001001110001000000011000100001111110000111111101010000000000000001010011001000000001010010000000100000000000000000000011000111000000000011010010000000000011010010001010110000000000011000110001011010101010011010010110001010010000000000000000000011010110101000000100000000001011011000000000000000000100000100000000010000000000101100110000000000000000000000011010001010011001000110011000110000000000101100100011011111011010110001001000010011110111100000011100000111100000010011110111100000110011110111001000010011111100100000110100110111100000111100000011011111111101000111100100111100000111100000111100100010010110011000000111100000000100100100010110110100000010011111011010110001100100111100000000010110110000000011011111010010110111110100111100000011011000111100000010010110011100100110100000101100000101100000111111111000000000000000000000000000111111111000000000111111111000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111000000000111111111111111111111111111000000000111111111000000000111111111111111111000000000000000000111111111000000000111111111111111111000000000000000000000000000000000000101100110110101100110100100000000000110100110000000000111100100000000000111110100000100000101100110101100100000000000111110100010100100111100110111110100110100110000000000011111001110110100000011111000000000111111110000000000000000010000000011101100100000000000100100100000000000000000000111000000111100010011000000111110100000000010100000010111111110100100100010000100000110010011011011011011001011011011000100001011001001001000011011011110100100000011011010000000011011011010011011010000000000011011011011011011011011011011010010011011001000000001001001001011011011111010010101101001001001011000100011000000000111000000011001011000000000001001011000000010000100011001001001011011011111011011001011011100100000111001011011011011011011011011011101011000000100111110000111010100111100011010001000111110011000001000111010000000000000101010111110100000111110000101010011010000000111100100111110100111110000111110100111110110100101000010110100111110100001110110000100000111010011010001011110001100100111100111110010000001100111000011010000011010001110101100100110110000001111000111110111000100000001110100111010000001110000010000011101010000000000000000001000000001001100110101111111101100010000000001001010010000000100101011111000000001000000000111101010000000001001000100000000100000000001000100000000110110111100000000000001000000000100111110000000001101100010001100010000000000000100001010000010100000011111101010111110010010000100000000111001000001000100001000000000000000100000000011000000000000000000100000000100100111000111111100101111100000000000101111000000000000101111000000000100101111000000000100101011100101111111010110000101111100101111100101111000101111100101111000000000100110111100101111000000001000001001100111111100000000111011001000000000100111111010010000000000011100000000100000100000101101100100011100000111101111111111000100000000001100100111100101011000100000100110010001011011011000000001011001101110111011001001100110000011011101100100000000011101111111111011011101001011001111110011011001101001001001001001000011011000001011001100110000000000000011011001001111111111111111011001001101110111101110111000111111001001001100111111111011111111110111101110111010000000001001011100011111011011001100110111001001111011001001000001001101101111000010000111111000111000001111000101000000000001000001000000000111000000000000000111001100000000000101000100101000100000000000111000000111010100101001000111000000001001100000000000111101000111000001000001000100000000111000000000001000000000000000000000111000101010000000000000000000010000000001000110110100010000000011111000111000100000010000001111000111010101111101100000000000110011101111111111011111011111011110111000001011111011110001101011111011100001111110011111011101001011111111111111111111101101011111011111111111011111111111111110111111111110001011011111111011111111101111110100001001111111001111000001111100101110100110111111011111111101111111011011001001111000001110011011011011011010010111111111111111101111111111111011111110110011111111111011010010110000000000010110100000000000000111111000000000010011100000000000010011111000000000010000100000000000000000000010011100000000000000000000000000000000000000000000000010011001000000000000000000111110110000001111001000000010010101010001111110010100011111110010011111010001000000011101000001111000000000000000000000000000000000000010110100010000110000000000000000000111101110000000000111111000011101000110101000001000010110001000000000000011111000000000100000011000011000000000011000011101000011000100011001000100101000100111000011111000111111000001000010000011000111101000000011001100000101111101000011000000101000010000000000111101000000000001100011000000000000101000100110111000111111000000101001011011000100000100000001100111101000100001000110100000000000000110110111100000011110100111000000000111101011000000000000000011000000000010100111000000000110100111010100111010000000100100111111100111111100111010000111111100111000000000001010111000100111000000000101101101100100111000000000001000000000000100100010111000000000100000110000000100010000000000111001111100111011000010100100111000100000011100000100100111010100111000000110000000110111111000111101000001111000000000001111000000000000110111001000000001111100111100000001000111111000110101000101000001111001000111111000101111000111001000101111000000000110111000000101001000001000000000111111101001000000000000000000100000001000111001000000000110011000000000000000000000111110100010111111000000111000111011000000000111000111010111001000100011000111000000000000000000001000000011001000001001000000000000001001000001000011001000000000000011101001000000000101001000011101001000000000001001001001101001111101001011001001001101001000000000001000000000001001100000000000000000001001001000000000000000000100000100000001001000000000000010000000000000000000000010010001000001000001001001001001001000000000011001000001000001011101001000000000000000000100111111000111001110111111111111101000011000000000000111111111010000100101111111111111111111111111110111111000000000111111111000000001000000000000011011111111111000000000110111111111111111111101111000000000111111111111111111000000000111111111111111111000000000000000000111111110111111101000001001111111111000000011111111111011000000000000011111111111000000011111111101000001000000110100110100000100110100000001000000000000001100000110110000001101010010110000000000000110100100010110000000000000100100100010100100010110100000100100010110100001001000011110111000100100000110110001001110110110100000000000000000000000110110110110100001101010000000000000000000000000000000000000000100100100010100000100100001111011100000000110110100110110000000000000010000000111001001111011001111001001010100100011000001010000000011001011010000000011001000000000000011001000011001001000000100111001001111001001111001001011001011111001000011000000011000000111001001111000000000000011011001001010100100000000100010000000111001001000000000000100000000100100010000100001001000001000000111011011111001001001000100111001111111000001111000000000000000000000000011011110011111111011011110001000000111111111001000000011111111000000000010011110000100010011011110011011110111100000011111110011011110011111110111111111011011110000000000001011000011011110000000010101000011011011110000000000001000000000000100011011111000000000111111010100000000001000001011011110001011110010111111011011111000000001011111111011011110001011110010011000000000100111110000100000000111111000000100111000000000000000100111111000000000000111110000000111111111111000011111000000000010111110000111110000011101000111111000111111000000100101101110000111110000011101011000000000011000000000000111000100000001110110011011000000000000000000000000100110000100011000000000111111000010110000011110000000100101011100000111110000111100000000000000000000000011010110111110010011100100000000000011110100000000000111110000000000000011110010000000100011110100011111110000000100011110000011010110111110110111110110011110010000000001011100110011110100011000011000000000111111100000000000000000000011101111011110010000100001011011100100000101000000000111100000111111110011111100111110010001001000011100010011110110011110010101000100111111111100110110111111110100110100111111111111110110111111111010110100111111111100110100111111111000110100000110100111111111110111100000110100000110100110111100000110100111111111010110110110110100111111101111111111111110110111111111111011011111111101111100110111111011111111110111111111111111111010111100000110110000101101100111100111111011111111111110111110000100100110110110111101100011111111011111011011111111010011000010111111111111111011111111011100110011111110111111100011111111011111111111111101011111010011111111011111111111111111011111111010110100000010111011111111111111110111011111011111111010011000111011110111111111011111111110111101111111111110101100110011100010011111001011111011111111011111111111111111111111111011111010011010111000011111010000010000111101101101000000111011010000000110110100010000010101111011010100010000111101000000000001111110000111111000000000111111001000111000010111111011111010000111011010000000011111001111111001000100111001010111111111100010000001100000000000100011111111001000000000110111000010000011010000000000000010000111111000011111011111001000000010000100111111111001000111001111011011010000000111001000101001100111001000000000000011001000000000000111011001000000010111011001001000110111111001111011001000000001111011000111001001111001001111011000111011000000000001110101000011001000000011001000010110011001000000000000000010010000010011011001000010000010001000010000000011000010010110001001111101000001011001011011001000010011000011001111001000111001001000000000000000000001001001001011011001001001000000000111011001000100100001001110000000000101001011000000100101001011101001001000000000001011010001011011001001001001011110001101001000000000000100001001101111001101000000000100101000111000000000000000000001001100101001011000000000001001001000000000000000000000001001101001000001111010001011110000000000011111100001000000101101010000000001100000011000000010010100001010011011010000000011001110100010100000001000100001110010110000111010111100000010000011110000001011000100110000100011111110000000110101110011110011110101100111111011010110101111010101110000101011001000110100011101101101111011110110100111111011010110101110110101001010110010111000011000011010101001110010100100100011010011010110100111110001010000101010001000010001100001011010001010111101001011000011010010100010001110100011110000111010100001111111110000101011010100110000101111111010000111000110110001110000101010111101010110111100111110101010010101111100111111111111011100110100101101111111110101010101000011111010111011000111101001110001101110000110010001010101010101010010011101001101100011110100100111101011000010100100110001011010010111110100011010100011011001101001111110000111011010000110011001001100010001010000110010111101110111011100111011111100110101011111110011010000111101111110010000111111111001000000101000100000000010010111010110101110001001100100100000000000101000110001010110101100011000001100000000010011000010000100000010000101000000101100000001010111010111111011101000100111101010010000010100100111010100110000111111011001110011010101101010100100100111001011010011000010001101110000110000110010111001111111010101101011111110110111101010110000010000100110110010010010110110111101011010101001100000000110110010010110100100100001001010001010000010001000110000100111101100011001011100100000010110000100000101001001011001010000001010001001110111010110111100111111010101101111111101110100011111110010111101001011111101110000011111101110110110100111001011010110101111001100000000010001111100001000111111111111111111101111100111001010010111110000100110110101010111110111111110011001100111110110110001101110101000110000101100101010101010100111010001111110111010000000010101110011101101101100101100011100111110100110100101001001110100110111110100011110000111111100010110100101011111001110000101101000001011010011111101001110101110001111111101110100001100011100100010110000010101010111100010110100001000001010001110011000110001000110011101000110110001000100010100000010010110111101111010001010010011100111101110001110011100110101000100101110100001010111101101111010001011010111010111101110011101010101110101100000101110110001100101111001101010001011010111110100101000011111001110110000010000110110100101011100001000110010000110111001110000000010011101000010010010000110010100100010000010000000000010000000000000110001100010001110000100000000100000100100000000011110000011111011011000100011100001000110000110001100010101100000101100001001011110110100111010011011010111111100101110100111111100111110001010101010110101010110010100111010001010001010110100001110000111010101110101000000101000000000011100001000110010000101010000110100001000011101000000100000000100010110100010010000001000010000000000001000010111101000000101001000100100100000001000100000110111100111011110111110001101101111000111010101011100010101111100111111001001000110110001111100010011011111110111101110001111110111110110111110111010110111010110000100001000001000000010010001000110000101000001010101100000100000000000010100001000110110000111011000110100000000001101000000100000000000010000100000111110010000011010010000010000110111100110100101001101101100100000001000100001110111111111111111011010111111111110101111010111111101110101111101111111001001011110100000111110010011011010110111101110101111111000100100101110101000100011101110101100010110010100100000110000000100000111001001010101100000100000000000101111001000101110000010110001110000000000011100100100111010110110010011111001100110011000101110011100110101111111101100011111001100101011100001100111100110010110010111111110101111011011110111101111000110111111100101101001101111100111011110111011001010011010101010110001010110101011001101011011100110110110000111001001011011100110100001100111110101001010010110100001111010110111010111101100100101000001010101110100001000001111010100000001010101001110111001101010001010101101111111100111110111101100001111011101100001111011111111111111000011011011011001111011100111110011101111001111011001101011100011101011111111111111011110011000100001100010100000101110101011010010101010100001000000100111010101010110000100001001000010100010010010000011010010001011010001000000101101000100000010010000000110010100010111001100001111011101000001010011001110111101001011101110111101110110010100010011011100101111011101101111011010001111101101001101000110011101001111010100000011001000101001010011001001001010000101101101001101000010011111111111110001100110001110110000000111101100100111011111111000110100001010011100001001101010001110010011100001110110101001110101000100000000101100100001011101101010010101010111001000011110001100000001011011101110111001001001001110101010110110010101010011101000111110011101101111011011001110101101001000000100001010000000010101010101101000001000000000100001011011001110100011000001000001100110110100011001111110010000011010000111110101011001110100000000101010110001110010111000110001011110010011010110101001010001001101100000010110101010101000110001010100101111111100000001000111011001110011000101101010111000110010101011100101011000001011111000010101100101011001011010001100111010100000110010111101100001010001101010111011111111100110101011111011000111111011111010011011111111111000011100100111110011111011101100101001111111100011101011101110000011111000101101001110010101110101101100001111010001111001101001001011111111010101011110110111100111011110111110000100001111011111010011000011010011111101110111101011101100011111011100101111010111100010111011110001100110010001001101110011110111001000000011110100010011111000100001111000101000000010001001101101000000110110001001001111000101110101101100011001011001100100011011001111111101010101001110111001001111000101110001101100001101011001111001110011001111111101011101011110101111111111100001011000111110010010101101101110111011111111010010100001111000111001111011100101010101100110011011010101110110111011101111111111010001011110111001011111000111110001100110101011010000110011110011001011011111010101011110011101010011100111100010110010100001110010111010110011111100000010010100010110010000101011111000000010100011010100100110101110011001110100000010101100110000001111001111000101100101011111010110111101101110110011101011111111000001110110001010001110010101010111101100010110001100001101010011101111101101001001010110100011001011000101010101001000010011010110011000011011010101110101010100001010110011011001110111111100010111101001111011111010000111111010011000111111111111101010110001100010011010110011100000111011111010100100111000010010111110100001001010101010010100000001011000010110101101101100010011100101100010000000110000001110001000010101000101101000010110001000000101011011001111101000001000100000101101010001000111110001101101101111011001111110111101111010111101010011111110101001010101100111110111011110111110101001111000100011101011110111010001111110101111011000010100110010000100011011000001011110011001001111111011011001111101001011011001110101010000111110111011100001101110111011101010110011000001010110011000000010010100010011101000011010000100001100110011000101101111000100000110011001101011010100000111101000011011010111001101010011000101111111001100000010001001001111010101100101100000011010010011100001000001011111110111010101001111001110011011101011001000010111101100010010111010110010011110010010000110010010111001111111110101110101111110101111111101111110110011111111111111011111111110111001110100010101010101101100111110101101111111111001101110111110011000011100111010000010010111010001101100001100001001100010011000111110111000010010010100100001010010000101111101011101000111111101010110111101111011011101011011111101110011111000110001101100010011110010101101111110010111110100011010110010110001001111001101101011011001001001111101110110011010011101011111111100000111011100000111000100001000001100010001111000100100100100010000011101011100101100110011000111000100011000001010010001010001100110000101010101010101101000101100100001000110001100011000001100010011010100101010000101010111110101101000101100101001000111000100111001101100010101101100101010010100100111111111111000101011111001101000001101101010111000001101110001110110011010001101000101101100110101000111010111001001111001111100010011011011100110010001110101010101010000111100011001010100101000111000001110010011010010100110000101110101000100000010101000000001110111101100111000001100010001010010100100000101010101010101010000101010101001100101111100101001001101011101010110101101010101101111110001011000111111111001100010110101101010111000100101101001110111111110001101010111010101010111011001110111010101111111111000110111101000011001111010101110111111110101111011111111001000001100100010010000110011100000111000101010100010101010000111010010110110110111011101101011111000100011101000100011010000101100011011010000110010111001001100001100100011011001110111011011100000110010111111001010001110110001010101111001111111011100011111101100101100111111011100011110110111111101011111111111110010110110100110001001011010001001111001111010000011110101101101011111110111001111000111011111111100001110001011010110110110111010010111011101110100011111100011010110110110111011011111101001111111111010010110111100111101010011111111001000010010110111100011011000011101101110101000011010101111101101101001010110001100100100101010001000011001111000101010001000001100100101100000001000101000000010000000001000001000000001010001100010001010011101010100000000100100100001000111001011101001001000010011010101100010001001000101110001001000101100001001010100101111101001001010010011010011100010010101110111010001011010110100001011001111000011100010011000110010110001010010110010101101001010011010010000111000010010110000001000001100100000011011100011001110000000011000101000101100010101110110110000011010101100110011011010100111001110001100010000101010101100010101111010010000001110011110100001011100101000100110001100100000100010100010100101101010011010000101010101101000111110001000100101111000000011101111101011001111101011010110001101011101100100101110001000110100101010001010111111101011011101110010110001001000001100100001011011100010000110001100010101101000101100010001010000010001101010001010010011101000110011101010100100110100101010100000110101011100011001111110011011111111110110110110111110100100101110111111111101110111011001100010010101010111101000011110011000011100111000100101101111001001010110101001100110010101110101101100001111011000011100011010101111111101010001111110110010100011001110001110100000011011110011001110101010000001101101101111010111011101111111001011011010100110101001010110001010101000010011000110110101011111011001010011100101110111101111011011011000011011110011101011011111010111111110011001101011010100100111101000011111000100100101110001001111101111001100010110011000100011010000110111101100011011000110000100110001001101101111001100000010101101100111010101010111101100011110001100100101111010101111111111001001011110111001100010010101110101101100011011000000101110111001001110111111011001010110000001101011000100100101101100010111000010100001000011001001000101001000010110101010101111101011001101101000000111000010000110010001110111000000101110010101001000011011100010111110110111000001110011101010100100110000001111110110010011011111100110010101000111101100011110011001001110000010111111111101001101011110001001111110110101110001101100001110011001111110111011101111111101011011111110111010100100000110110001111100101101000100110010101000111110111111011010110111110011110100010110110101010101000110111101110010001100110100001001001011110111110010110100011111011110111011001010110101011010001100110010001000101011110101000001110000101010111110001111010010010000011010001110110001100100110100100001100100011000101000100110010111000110110010011001000100110000100000101110100001010110101000111000101111010101010110101101001001000100110100011000101011100001110011110000011000001111011101000110111101011000001110110000100001101011110111100010010000100110100101011100010101111001011010001110100001100101001111100110100101100000101011111110000010011010010000010000001100010010110000011000101001100010111000101010001100110011010010100010000101001100100000000000101010100001110111111100111000001110110001010110100100110101011101110100001000101010110001110010101100010100000110011000010110101100000101011001100100101010001000010000111010100100010100010111101000011011000100000101011001000101101000001000000000100111010001001011111100000111000010010010010010000100010000010000110110110001100011100001101011111100010111010110110110111100101100110100010000111010111001100101010101101001011000110111100000100100101000100100111010010010110010111001011001110000000101110101101100011111010100100100111011001010101011000000011100101001000011001111011100100101101001010010101010001000011011110101000000011110010011111010101010101110000101000010010110010100001000010001000000110100000001110111110101101011111100110111100001010011010000101110010100010010110111011011001101010001101010111000110111101000110000111010100100111010000110110011110001000011100001001001110100100110101000000000110000000010010010010010110100011000110001110100101011111010010111101010000000010000100110111010010000111011111001000101111000001000110101000010010010010000010000001100010000000010001100000001010101101111101011001111001110011010010011011111000110010001010111111111011010011001111011100111110111101111101111111010111110110011101011111111010111011110101011110010010111110001001100111111111001010100001010101110111101011011111100110001100000010100110101011100011110111000101100011010000100001100101001110111001011010000101011110111100110011000111000101000100110011011101110011100111010001101001011110111011110100110011000110000111100110000001010111110011101011100101000001011110110010111100000011011100100101111111000001000101010000000000100010010100011010011010011101000010010000100100111111000000100101010001000000000100111000110011011010111100000010001010100010100101000000001101000000000000000011011100111100111010111100110011010011000101000100010001001111111000001011110011011101111110111110111101101111111011010111110111010101111111111011111011110001011011111010111110011101100001101111001111010101010111111111101011101010110101101010111100111110001111111101101011011111010101110111010110101010111011111100100110000111111011111110111101101111000111110001110111010111011111010110111001010010010000110010110111100011111111000101100011010001010101101011000111110100010000100010100010101001000011101101000001101011100101110101001001010100101010110101110011000001111011000010110101100000101010001100101101000101100100001110111010111101001101100001101111010000110010001100101010001010000110111111011111101100101101111111110110111011010110100111110110110111110011110111010111011010110010000001110000101111010010100111000001100001110100000101001001011110111100110010000010100001100010001010111101100010100011111100100001001001011101101110110010000011010011010010000011100100100000010001100111110000000101010100001110111010100101111001011111101001100111101010100001100110001111101111011111111000111100010011100101011011100011110111100001101011011100001111101011101110111000110000000001010011110100010010000100000001000100100001000001010011010100001100010010000001010001100010000010100100110000111011100010100000000101000100001110111111101111001001110010111010010101111010101010101110100001000101110101001010110100100111010001110010011010111101110000101010110100100001010101000110001010110100000011010001010001000010110000100000100011001000100001000101000000001010011011110110101100011010111100101101011111111110011101111000001010010010110001000000100010001100000001001110101101011000001010001011111000001000010101000111001111000000101111000010101101000000001111011010111111111010001010011111110101011110110100101110000100110101000010001011001100011001110011111010011011110011001101111010101100001000011101001100001100101110011001110010101000011011110001111011100111001101000110011100101100011100101110001111111000010110100011011100100110101101011101000110111100000010011110010100001010001010010110101001011101000100001100001100000010110001000000010111000100011000010010010110111111010000000101100000001100001001100000000000001010001000010001010010010000001001010101001010001100001100000110111001000000011111100000011011011010001010011111000011001011110110101100001011111100101110111100111110011001011010111010001010110011000101111100011100011101110000001010101100011110011010001000111100100000010101000100111101011101000100110101001010011111010100100011011010111110100001110111001011000000110010011100100100100011101111011110010001010010010010011101110110011011110000101100101011001100100011101010101010011000001011101010011101111000110101000011001101010011011100101101111100111010001011110000000010110000101100111011100101001101000010101100001100101110001001101011011010000110110101001100000010101101110101000010111100000111011110010100110110011010001010011100110001001101000000000100110001110010001000100001001110011001010110110000000001010011010001011011000000000101000101001000110001110110001011101000010000100001000000100010011011001101010010011100001100111100111010101010100010011100011011111000001001011101001101000010011000001100011100000100111010001000010100101001001001001000001100011100100100110000000000011111010100010001010010010010000001000101001011001001001010000100110100000000001110000100000011010010010010010101000100110011101101000000000010111100101110111111111110001111010000010010110110000011010100111100111110011011101100100111010110011100110101000001101010011000111110010110110000111000011111100100100101100000010001110000101001101000010000110101011100101000101111000101100101000001101110000101000001010010111010011011011101001000001110101110000101100001000000001110101111000001110011011010000011100010000001111010000010011101000100001000111100011011100000101001111010100000010110110110000001001001010010001101000101111110001011100111010011010111110001101100101110100001001101000000001111100011001010000010100111010010000010011101001100001110100000101100101001101101001011001111000010011101000111111010011111110001010010011000110100001001110100001010011101010000010101010110111010001001110011000001011110010010000010010111001010110101011100000001010000110000110000000100111110101101001101000010111100001010011110000100100010001000000110111000011011101111011101001101000110111000000000010010000100111010000010111110111011010101001101011000101010010100110000000001010111011100010001010010111010100001110101011010001001111110010110101100101111111111010001100111010111101010011101101110010011001101010101010010111100100111011111010000110111000001000001111100111011100001001101001000011011100101000110110000001100100000101000111100100000010011000101111100000000111101110010000011010100001110011011011011111010101000110001001100110010101100111001000011111001000000001110011001011100111010101011010000110010111111000101010010011110001101111011011110111110001011000011111111001010010110001111010001010010001100001100110001111001110110100001010100000000001011010100011101001010010010000100000101100100001100100101010000110100000000101000010100010010000001011101000110100001100000001011001001110001100001000000001000110101100011000101001011000010110101100000101011101110100000000101010000001010110101100111000001110011001011100101110000101010110110101000000101100000011011110000101101001001010000011100000000010010001111100011001010010110000000001";

begin

top_inst: entity work.top
    port map (
        clk         => clk,
        reset       => reset,

        w_en        => w_en,
        w_in        => w_in,
        w_out       => w_out,

        row_in      => row_in,
        ready       => ready,

        row_out     => row_out,
        done        => done
    );

    clk   <= not clk after CLK_PERIOD/2;

    -- Load weights
    process
    begin
        w_en <= '0';
        w_in <= '0';

        wait for 2*CLK_PERIOD; --reset

        for I in 0 to WEIGHTS'length-1 loop
            w_en <= '1';
            w_in <= WEIGHTS(I);
            wait for CLK_PERIOD;
        end loop;
        w_en <= '0';

        wait;
    end process;

end architecture;
